module RISCV_Single_Cycle(
    input         clk,
    input         rst_n
);
// Đây là module top, bạn sẽ tự kết nối các module nhỏ ở trên theo sơ đồ single-cycle CPU.
// Do mỗi lab, mỗi thầy sẽ có sơ đồ và tín hiệu riêng, dưới đây chỉ là ví dụ tối giản.
endmodule
